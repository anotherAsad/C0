/* VERY VERY BRAIN-UNFRIENDLY CODE FOLLOWS */
module instrMUX(out,
	i00, i01, i02, i03, i04, i05, i06, i07, i08, i09, i0A, i0B, i0C, i0D, i0E, i0F,
	i10, i11, i12, i13, i14, i15, i16, i17, i18, i19, i1A, i1B, i1C, i1D, i1E, i1F,
	i20, i21, i22, i23, i24, i25, i26, i27, i28, i29, i2A, i2B, i2C, i2D, i2E, i2F,
	i30, i31, i32, i33, i34, i35, i36, i37, i38, i39, i3A, i3B, i3C, i3D, i3E, i3F,
	i40, i41, i42, i43, i44, i45, i46, i47, i48, i49, i4A, i4B, i4C, i4D, i4E, i4F,
	i50, i51, i52, i53, i54, i55, i56, i57, i58, i59, i5A, i5B, i5C, i5D, i5E, i5F,
	i60, i61, i62, i63, i64, i65, i66, i67, i68, i69, i6A, i6B, i6C, i6D, i6E, i6F,
	i70, i71, i72, i73, i74, i75, i76, i77, i78, i79, i7A, i7B, i7C, i7D, i7E, i7F,
	i80, i81, i82, i83, i84, i85, i86, i87, i88, i89, i8A, i8B, i8C, i8D, i8E, i8F,
	i90, i91, i92, i93, i94, i95, i96, i97, i98, i99, i9A, i9B, i9C, i9D, i9E, i9F,
	iA0, iA1, iA2, iA3, iA4, iA5, iA6, iA7, iA8, iA9, iAA, iAB, iAC, iAD, iAE, iAF,
	iB0, iB1, iB2, iB3, iB4, iB5, iB6, iB7, iB8, iB9, iBA, iBB, iBC, iBD, iBE, iBF,
	iC0, iC1, iC2, iC3, iC4, iC5, iC6, iC7, iC8, iC9, iCA, iCB, iCC, iCD, iCE, iCF,
	iD0, iD1, iD2, iD3, iD4, iD5, iD6, iD7, iD8, iD9, iDA, iDB, iDC, iDD, iDE, iDF,
	iE0, iE1, iE2, iE3, iE4, iE5, iE6, iE7, iE8, iE9, iEA, iEB, iEC, iED, iEE, iEF,
	iF0, iF1, iF2, iF3, iF4, iF5, iF6, iF7, iF8, iF9, iFA, iFB, iFC, iFD, iFE, iFF,
	S);
	output [20:0] out;
	input  [20:0] i00, i01, i02, i03, i04, i05, i06, i07, i08, i09, i0A, i0B, i0C, i0D, i0E, i0F,
				  i10, i11, i12, i13, i14, i15, i16, i17, i18, i19, i1A, i1B, i1C, i1D, i1E, i1F,
				  i20, i21, i22, i23, i24, i25, i26, i27, i28, i29, i2A, i2B, i2C, i2D, i2E, i2F,
				  i30, i31, i32, i33, i34, i35, i36, i37, i38, i39, i3A, i3B, i3C, i3D, i3E, i3F,
				  i40, i41, i42, i43, i44, i45, i46, i47, i48, i49, i4A, i4B, i4C, i4D, i4E, i4F,
				  i50, i51, i52, i53, i54, i55, i56, i57, i58, i59, i5A, i5B, i5C, i5D, i5E, i5F,
				  i60, i61, i62, i63, i64, i65, i66, i67, i68, i69, i6A, i6B, i6C, i6D, i6E, i6F,
				  i70, i71, i72, i73, i74, i75, i76, i77, i78, i79, i7A, i7B, i7C, i7D, i7E, i7F,
				  i80, i81, i82, i83, i84, i85, i86, i87, i88, i89, i8A, i8B, i8C, i8D, i8E, i8F,
				  i90, i91, i92, i93, i94, i95, i96, i97, i98, i99, i9A, i9B, i9C, i9D, i9E, i9F,
				  iA0, iA1, iA2, iA3, iA4, iA5, iA6, iA7, iA8, iA9, iAA, iAB, iAC, iAD, iAE, iAF,
				  iB0, iB1, iB2, iB3, iB4, iB5, iB6, iB7, iB8, iB9, iBA, iBB, iBC, iBD, iBE, iBF,
				  iC0, iC1, iC2, iC3, iC4, iC5, iC6, iC7, iC8, iC9, iCA, iCB, iCC, iCD, iCE, iCF,
				  iD0, iD1, iD2, iD3, iD4, iD5, iD6, iD7, iD8, iD9, iDA, iDB, iDC, iDD, iDE, iDF,
				  iE0, iE1, iE2, iE3, iE4, iE5, iE6, iE7, iE8, iE9, iEA, iEB, iEC, iED, iEE, iEF,
				  iF0, iF1, iF2, iF3, iF4, iF5, iF6, iF7, iF8, iF9, iFA, iFB, iFC, iFD, iFE, iFF;
	input  [7:0]  S;

bitmux256 MX0(out[0], {i00[0], i01[0], i02[0], i03[0], i04[0], i05[0], i06[0], i07[0],
i08[0], i09[0], i0A[0], i0B[0], i0C[0], i0D[0], i0E[0], i0F[0],
i10[0], i11[0], i12[0], i13[0], i14[0], i15[0], i16[0], i17[0],
i18[0], i19[0], i1A[0], i1B[0], i1C[0], i1D[0], i1E[0], i1F[0],
i20[0], i21[0], i22[0], i23[0], i24[0], i25[0], i26[0], i27[0],
i28[0], i29[0], i2A[0], i2B[0], i2C[0], i2D[0], i2E[0], i2F[0],
i30[0], i31[0], i32[0], i33[0], i34[0], i35[0], i36[0], i37[0],
i38[0], i39[0], i3A[0], i3B[0], i3C[0], i3D[0], i3E[0], i3F[0],
i40[0], i41[0], i42[0], i43[0], i44[0], i45[0], i46[0], i47[0],
i48[0], i49[0], i4A[0], i4B[0], i4C[0], i4D[0], i4E[0], i4F[0],
i50[0], i51[0], i52[0], i53[0], i54[0], i55[0], i56[0], i57[0],
i58[0], i59[0], i5A[0], i5B[0], i5C[0], i5D[0], i5E[0], i5F[0],
i60[0], i61[0], i62[0], i63[0], i64[0], i65[0], i66[0], i67[0],
i68[0], i69[0], i6A[0], i6B[0], i6C[0], i6D[0], i6E[0], i6F[0],
i70[0], i71[0], i72[0], i73[0], i74[0], i75[0], i76[0], i77[0],
i78[0], i79[0], i7A[0], i7B[0], i7C[0], i7D[0], i7E[0], i7F[0],
i80[0], i81[0], i82[0], i83[0], i84[0], i85[0], i86[0], i87[0],
i88[0], i89[0], i8A[0], i8B[0], i8C[0], i8D[0], i8E[0], i8F[0],
i90[0], i91[0], i92[0], i93[0], i94[0], i95[0], i96[0], i97[0],
i98[0], i99[0], i9A[0], i9B[0], i9C[0], i9D[0], i9E[0], i9F[0],
iA0[0], iA1[0], iA2[0], iA3[0], iA4[0], iA5[0], iA6[0], iA7[0],
iA8[0], iA9[0], iAA[0], iAB[0], iAC[0], iAD[0], iAE[0], iAF[0],
iB0[0], iB1[0], iB2[0], iB3[0], iB4[0], iB5[0], iB6[0], iB7[0],
iB8[0], iB9[0], iBA[0], iBB[0], iBC[0], iBD[0], iBE[0], iBF[0],
iC0[0], iC1[0], iC2[0], iC3[0], iC4[0], iC5[0], iC6[0], iC7[0],
iC8[0], iC9[0], iCA[0], iCB[0], iCC[0], iCD[0], iCE[0], iCF[0],
iD0[0], iD1[0], iD2[0], iD3[0], iD4[0], iD5[0], iD6[0], iD7[0],
iD8[0], iD9[0], iDA[0], iDB[0], iDC[0], iDD[0], iDE[0], iDF[0],
iE0[0], iE1[0], iE2[0], iE3[0], iE4[0], iE5[0], iE6[0], iE7[0],
iE8[0], iE9[0], iEA[0], iEB[0], iEC[0], iED[0], iEE[0], iEF[0],
iF0[0], iF1[0], iF2[0], iF3[0], iF4[0], iF5[0], iF6[0], iF7[0],
iF8[0], iF9[0], iFA[0], iFB[0], iFC[0], iFD[0], iFE[0], iFF[0]}, S);


bitmux256 MX1(out[1], {
i00[1], i01[1], i02[1], i03[1], i04[1], i05[1], i06[1], i07[1],
i08[1], i09[1], i0A[1], i0B[1], i0C[1], i0D[1], i0E[1], i0F[1],
i10[1], i11[1], i12[1], i13[1], i14[1], i15[1], i16[1], i17[1],
i18[1], i19[1], i1A[1], i1B[1], i1C[1], i1D[1], i1E[1], i1F[1],
i20[1], i21[1], i22[1], i23[1], i24[1], i25[1], i26[1], i27[1],
i28[1], i29[1], i2A[1], i2B[1], i2C[1], i2D[1], i2E[1], i2F[1],
i30[1], i31[1], i32[1], i33[1], i34[1], i35[1], i36[1], i37[1],
i38[1], i39[1], i3A[1], i3B[1], i3C[1], i3D[1], i3E[1], i3F[1],
i40[1], i41[1], i42[1], i43[1], i44[1], i45[1], i46[1], i47[1],
i48[1], i49[1], i4A[1], i4B[1], i4C[1], i4D[1], i4E[1], i4F[1],
i50[1], i51[1], i52[1], i53[1], i54[1], i55[1], i56[1], i57[1],
i58[1], i59[1], i5A[1], i5B[1], i5C[1], i5D[1], i5E[1], i5F[1],
i60[1], i61[1], i62[1], i63[1], i64[1], i65[1], i66[1], i67[1],
i68[1], i69[1], i6A[1], i6B[1], i6C[1], i6D[1], i6E[1], i6F[1],
i70[1], i71[1], i72[1], i73[1], i74[1], i75[1], i76[1], i77[1],
i78[1], i79[1], i7A[1], i7B[1], i7C[1], i7D[1], i7E[1], i7F[1],
i80[1], i81[1], i82[1], i83[1], i84[1], i85[1], i86[1], i87[1],
i88[1], i89[1], i8A[1], i8B[1], i8C[1], i8D[1], i8E[1], i8F[1],
i90[1], i91[1], i92[1], i93[1], i94[1], i95[1], i96[1], i97[1],
i98[1], i99[1], i9A[1], i9B[1], i9C[1], i9D[1], i9E[1], i9F[1],
iA0[1], iA1[1], iA2[1], iA3[1], iA4[1], iA5[1], iA6[1], iA7[1],
iA8[1], iA9[1], iAA[1], iAB[1], iAC[1], iAD[1], iAE[1], iAF[1],
iB0[1], iB1[1], iB2[1], iB3[1], iB4[1], iB5[1], iB6[1], iB7[1],
iB8[1], iB9[1], iBA[1], iBB[1], iBC[1], iBD[1], iBE[1], iBF[1],
iC0[1], iC1[1], iC2[1], iC3[1], iC4[1], iC5[1], iC6[1], iC7[1],
iC8[1], iC9[1], iCA[1], iCB[1], iCC[1], iCD[1], iCE[1], iCF[1],
iD0[1], iD1[1], iD2[1], iD3[1], iD4[1], iD5[1], iD6[1], iD7[1],
iD8[1], iD9[1], iDA[1], iDB[1], iDC[1], iDD[1], iDE[1], iDF[1],
iE0[1], iE1[1], iE2[1], iE3[1], iE4[1], iE5[1], iE6[1], iE7[1],
iE8[1], iE9[1], iEA[1], iEB[1], iEC[1], iED[1], iEE[1], iEF[1],
iF0[1], iF1[1], iF2[1], iF3[1], iF4[1], iF5[1], iF6[1], iF7[1],
iF8[1], iF9[1], iFA[1], iFB[1], iFC[1], iFD[1], iFE[1], iFF[1]
}, S);


bitmux256 MX2(out[2], {
i00[2], i01[2], i02[2], i03[2], i04[2], i05[2], i06[2], i07[2],
i08[2], i09[2], i0A[2], i0B[2], i0C[2], i0D[2], i0E[2], i0F[2],
i10[2], i11[2], i12[2], i13[2], i14[2], i15[2], i16[2], i17[2],
i18[2], i19[2], i1A[2], i1B[2], i1C[2], i1D[2], i1E[2], i1F[2],
i20[2], i21[2], i22[2], i23[2], i24[2], i25[2], i26[2], i27[2],
i28[2], i29[2], i2A[2], i2B[2], i2C[2], i2D[2], i2E[2], i2F[2],
i30[2], i31[2], i32[2], i33[2], i34[2], i35[2], i36[2], i37[2],
i38[2], i39[2], i3A[2], i3B[2], i3C[2], i3D[2], i3E[2], i3F[2],
i40[2], i41[2], i42[2], i43[2], i44[2], i45[2], i46[2], i47[2],
i48[2], i49[2], i4A[2], i4B[2], i4C[2], i4D[2], i4E[2], i4F[2],
i50[2], i51[2], i52[2], i53[2], i54[2], i55[2], i56[2], i57[2],
i58[2], i59[2], i5A[2], i5B[2], i5C[2], i5D[2], i5E[2], i5F[2],
i60[2], i61[2], i62[2], i63[2], i64[2], i65[2], i66[2], i67[2],
i68[2], i69[2], i6A[2], i6B[2], i6C[2], i6D[2], i6E[2], i6F[2],
i70[2], i71[2], i72[2], i73[2], i74[2], i75[2], i76[2], i77[2],
i78[2], i79[2], i7A[2], i7B[2], i7C[2], i7D[2], i7E[2], i7F[2],
i80[2], i81[2], i82[2], i83[2], i84[2], i85[2], i86[2], i87[2],
i88[2], i89[2], i8A[2], i8B[2], i8C[2], i8D[2], i8E[2], i8F[2],
i90[2], i91[2], i92[2], i93[2], i94[2], i95[2], i96[2], i97[2],
i98[2], i99[2], i9A[2], i9B[2], i9C[2], i9D[2], i9E[2], i9F[2],
iA0[2], iA1[2], iA2[2], iA3[2], iA4[2], iA5[2], iA6[2], iA7[2],
iA8[2], iA9[2], iAA[2], iAB[2], iAC[2], iAD[2], iAE[2], iAF[2],
iB0[2], iB1[2], iB2[2], iB3[2], iB4[2], iB5[2], iB6[2], iB7[2],
iB8[2], iB9[2], iBA[2], iBB[2], iBC[2], iBD[2], iBE[2], iBF[2],
iC0[2], iC1[2], iC2[2], iC3[2], iC4[2], iC5[2], iC6[2], iC7[2],
iC8[2], iC9[2], iCA[2], iCB[2], iCC[2], iCD[2], iCE[2], iCF[2],
iD0[2], iD1[2], iD2[2], iD3[2], iD4[2], iD5[2], iD6[2], iD7[2],
iD8[2], iD9[2], iDA[2], iDB[2], iDC[2], iDD[2], iDE[2], iDF[2],
iE0[2], iE1[2], iE2[2], iE3[2], iE4[2], iE5[2], iE6[2], iE7[2],
iE8[2], iE9[2], iEA[2], iEB[2], iEC[2], iED[2], iEE[2], iEF[2],
iF0[2], iF1[2], iF2[2], iF3[2], iF4[2], iF5[2], iF6[2], iF7[2],
iF8[2], iF9[2], iFA[2], iFB[2], iFC[2], iFD[2], iFE[2], iFF[2]
}, S);


bitmux256 MX3(out[3], {
i00[3], i01[3], i02[3], i03[3], i04[3], i05[3], i06[3], i07[3],
i08[3], i09[3], i0A[3], i0B[3], i0C[3], i0D[3], i0E[3], i0F[3],
i10[3], i11[3], i12[3], i13[3], i14[3], i15[3], i16[3], i17[3],
i18[3], i19[3], i1A[3], i1B[3], i1C[3], i1D[3], i1E[3], i1F[3],
i20[3], i21[3], i22[3], i23[3], i24[3], i25[3], i26[3], i27[3],
i28[3], i29[3], i2A[3], i2B[3], i2C[3], i2D[3], i2E[3], i2F[3],
i30[3], i31[3], i32[3], i33[3], i34[3], i35[3], i36[3], i37[3],
i38[3], i39[3], i3A[3], i3B[3], i3C[3], i3D[3], i3E[3], i3F[3],
i40[3], i41[3], i42[3], i43[3], i44[3], i45[3], i46[3], i47[3],
i48[3], i49[3], i4A[3], i4B[3], i4C[3], i4D[3], i4E[3], i4F[3],
i50[3], i51[3], i52[3], i53[3], i54[3], i55[3], i56[3], i57[3],
i58[3], i59[3], i5A[3], i5B[3], i5C[3], i5D[3], i5E[3], i5F[3],
i60[3], i61[3], i62[3], i63[3], i64[3], i65[3], i66[3], i67[3],
i68[3], i69[3], i6A[3], i6B[3], i6C[3], i6D[3], i6E[3], i6F[3],
i70[3], i71[3], i72[3], i73[3], i74[3], i75[3], i76[3], i77[3],
i78[3], i79[3], i7A[3], i7B[3], i7C[3], i7D[3], i7E[3], i7F[3],
i80[3], i81[3], i82[3], i83[3], i84[3], i85[3], i86[3], i87[3],
i88[3], i89[3], i8A[3], i8B[3], i8C[3], i8D[3], i8E[3], i8F[3],
i90[3], i91[3], i92[3], i93[3], i94[3], i95[3], i96[3], i97[3],
i98[3], i99[3], i9A[3], i9B[3], i9C[3], i9D[3], i9E[3], i9F[3],
iA0[3], iA1[3], iA2[3], iA3[3], iA4[3], iA5[3], iA6[3], iA7[3],
iA8[3], iA9[3], iAA[3], iAB[3], iAC[3], iAD[3], iAE[3], iAF[3],
iB0[3], iB1[3], iB2[3], iB3[3], iB4[3], iB5[3], iB6[3], iB7[3],
iB8[3], iB9[3], iBA[3], iBB[3], iBC[3], iBD[3], iBE[3], iBF[3],
iC0[3], iC1[3], iC2[3], iC3[3], iC4[3], iC5[3], iC6[3], iC7[3],
iC8[3], iC9[3], iCA[3], iCB[3], iCC[3], iCD[3], iCE[3], iCF[3],
iD0[3], iD1[3], iD2[3], iD3[3], iD4[3], iD5[3], iD6[3], iD7[3],
iD8[3], iD9[3], iDA[3], iDB[3], iDC[3], iDD[3], iDE[3], iDF[3],
iE0[3], iE1[3], iE2[3], iE3[3], iE4[3], iE5[3], iE6[3], iE7[3],
iE8[3], iE9[3], iEA[3], iEB[3], iEC[3], iED[3], iEE[3], iEF[3],
iF0[3], iF1[3], iF2[3], iF3[3], iF4[3], iF5[3], iF6[3], iF7[3],
iF8[3], iF9[3], iFA[3], iFB[3], iFC[3], iFD[3], iFE[3], iFF[3]
}, S);


bitmux256 MX4(out[4], {
i00[4], i01[4], i02[4], i03[4], i04[4], i05[4], i06[4], i07[4],
i08[4], i09[4], i0A[4], i0B[4], i0C[4], i0D[4], i0E[4], i0F[4],
i10[4], i11[4], i12[4], i13[4], i14[4], i15[4], i16[4], i17[4],
i18[4], i19[4], i1A[4], i1B[4], i1C[4], i1D[4], i1E[4], i1F[4],
i20[4], i21[4], i22[4], i23[4], i24[4], i25[4], i26[4], i27[4],
i28[4], i29[4], i2A[4], i2B[4], i2C[4], i2D[4], i2E[4], i2F[4],
i30[4], i31[4], i32[4], i33[4], i34[4], i35[4], i36[4], i37[4],
i38[4], i39[4], i3A[4], i3B[4], i3C[4], i3D[4], i3E[4], i3F[4],
i40[4], i41[4], i42[4], i43[4], i44[4], i45[4], i46[4], i47[4],
i48[4], i49[4], i4A[4], i4B[4], i4C[4], i4D[4], i4E[4], i4F[4],
i50[4], i51[4], i52[4], i53[4], i54[4], i55[4], i56[4], i57[4],
i58[4], i59[4], i5A[4], i5B[4], i5C[4], i5D[4], i5E[4], i5F[4],
i60[4], i61[4], i62[4], i63[4], i64[4], i65[4], i66[4], i67[4],
i68[4], i69[4], i6A[4], i6B[4], i6C[4], i6D[4], i6E[4], i6F[4],
i70[4], i71[4], i72[4], i73[4], i74[4], i75[4], i76[4], i77[4],
i78[4], i79[4], i7A[4], i7B[4], i7C[4], i7D[4], i7E[4], i7F[4],
i80[4], i81[4], i82[4], i83[4], i84[4], i85[4], i86[4], i87[4],
i88[4], i89[4], i8A[4], i8B[4], i8C[4], i8D[4], i8E[4], i8F[4],
i90[4], i91[4], i92[4], i93[4], i94[4], i95[4], i96[4], i97[4],
i98[4], i99[4], i9A[4], i9B[4], i9C[4], i9D[4], i9E[4], i9F[4],
iA0[4], iA1[4], iA2[4], iA3[4], iA4[4], iA5[4], iA6[4], iA7[4],
iA8[4], iA9[4], iAA[4], iAB[4], iAC[4], iAD[4], iAE[4], iAF[4],
iB0[4], iB1[4], iB2[4], iB3[4], iB4[4], iB5[4], iB6[4], iB7[4],
iB8[4], iB9[4], iBA[4], iBB[4], iBC[4], iBD[4], iBE[4], iBF[4],
iC0[4], iC1[4], iC2[4], iC3[4], iC4[4], iC5[4], iC6[4], iC7[4],
iC8[4], iC9[4], iCA[4], iCB[4], iCC[4], iCD[4], iCE[4], iCF[4],
iD0[4], iD1[4], iD2[4], iD3[4], iD4[4], iD5[4], iD6[4], iD7[4],
iD8[4], iD9[4], iDA[4], iDB[4], iDC[4], iDD[4], iDE[4], iDF[4],
iE0[4], iE1[4], iE2[4], iE3[4], iE4[4], iE5[4], iE6[4], iE7[4],
iE8[4], iE9[4], iEA[4], iEB[4], iEC[4], iED[4], iEE[4], iEF[4],
iF0[4], iF1[4], iF2[4], iF3[4], iF4[4], iF5[4], iF6[4], iF7[4],
iF8[4], iF9[4], iFA[4], iFB[4], iFC[4], iFD[4], iFE[4], iFF[4]
}, S);


bitmux256 MX5(out[5], {
i00[5], i01[5], i02[5], i03[5], i04[5], i05[5], i06[5], i07[5],
i08[5], i09[5], i0A[5], i0B[5], i0C[5], i0D[5], i0E[5], i0F[5],
i10[5], i11[5], i12[5], i13[5], i14[5], i15[5], i16[5], i17[5],
i18[5], i19[5], i1A[5], i1B[5], i1C[5], i1D[5], i1E[5], i1F[5],
i20[5], i21[5], i22[5], i23[5], i24[5], i25[5], i26[5], i27[5],
i28[5], i29[5], i2A[5], i2B[5], i2C[5], i2D[5], i2E[5], i2F[5],
i30[5], i31[5], i32[5], i33[5], i34[5], i35[5], i36[5], i37[5],
i38[5], i39[5], i3A[5], i3B[5], i3C[5], i3D[5], i3E[5], i3F[5],
i40[5], i41[5], i42[5], i43[5], i44[5], i45[5], i46[5], i47[5],
i48[5], i49[5], i4A[5], i4B[5], i4C[5], i4D[5], i4E[5], i4F[5],
i50[5], i51[5], i52[5], i53[5], i54[5], i55[5], i56[5], i57[5],
i58[5], i59[5], i5A[5], i5B[5], i5C[5], i5D[5], i5E[5], i5F[5],
i60[5], i61[5], i62[5], i63[5], i64[5], i65[5], i66[5], i67[5],
i68[5], i69[5], i6A[5], i6B[5], i6C[5], i6D[5], i6E[5], i6F[5],
i70[5], i71[5], i72[5], i73[5], i74[5], i75[5], i76[5], i77[5],
i78[5], i79[5], i7A[5], i7B[5], i7C[5], i7D[5], i7E[5], i7F[5],
i80[5], i81[5], i82[5], i83[5], i84[5], i85[5], i86[5], i87[5],
i88[5], i89[5], i8A[5], i8B[5], i8C[5], i8D[5], i8E[5], i8F[5],
i90[5], i91[5], i92[5], i93[5], i94[5], i95[5], i96[5], i97[5],
i98[5], i99[5], i9A[5], i9B[5], i9C[5], i9D[5], i9E[5], i9F[5],
iA0[5], iA1[5], iA2[5], iA3[5], iA4[5], iA5[5], iA6[5], iA7[5],
iA8[5], iA9[5], iAA[5], iAB[5], iAC[5], iAD[5], iAE[5], iAF[5],
iB0[5], iB1[5], iB2[5], iB3[5], iB4[5], iB5[5], iB6[5], iB7[5],
iB8[5], iB9[5], iBA[5], iBB[5], iBC[5], iBD[5], iBE[5], iBF[5],
iC0[5], iC1[5], iC2[5], iC3[5], iC4[5], iC5[5], iC6[5], iC7[5],
iC8[5], iC9[5], iCA[5], iCB[5], iCC[5], iCD[5], iCE[5], iCF[5],
iD0[5], iD1[5], iD2[5], iD3[5], iD4[5], iD5[5], iD6[5], iD7[5],
iD8[5], iD9[5], iDA[5], iDB[5], iDC[5], iDD[5], iDE[5], iDF[5],
iE0[5], iE1[5], iE2[5], iE3[5], iE4[5], iE5[5], iE6[5], iE7[5],
iE8[5], iE9[5], iEA[5], iEB[5], iEC[5], iED[5], iEE[5], iEF[5],
iF0[5], iF1[5], iF2[5], iF3[5], iF4[5], iF5[5], iF6[5], iF7[5],
iF8[5], iF9[5], iFA[5], iFB[5], iFC[5], iFD[5], iFE[5], iFF[5]
}, S);


bitmux256 MX6(out[6], {
i00[6], i01[6], i02[6], i03[6], i04[6], i05[6], i06[6], i07[6],
i08[6], i09[6], i0A[6], i0B[6], i0C[6], i0D[6], i0E[6], i0F[6],
i10[6], i11[6], i12[6], i13[6], i14[6], i15[6], i16[6], i17[6],
i18[6], i19[6], i1A[6], i1B[6], i1C[6], i1D[6], i1E[6], i1F[6],
i20[6], i21[6], i22[6], i23[6], i24[6], i25[6], i26[6], i27[6],
i28[6], i29[6], i2A[6], i2B[6], i2C[6], i2D[6], i2E[6], i2F[6],
i30[6], i31[6], i32[6], i33[6], i34[6], i35[6], i36[6], i37[6],
i38[6], i39[6], i3A[6], i3B[6], i3C[6], i3D[6], i3E[6], i3F[6],
i40[6], i41[6], i42[6], i43[6], i44[6], i45[6], i46[6], i47[6],
i48[6], i49[6], i4A[6], i4B[6], i4C[6], i4D[6], i4E[6], i4F[6],
i50[6], i51[6], i52[6], i53[6], i54[6], i55[6], i56[6], i57[6],
i58[6], i59[6], i5A[6], i5B[6], i5C[6], i5D[6], i5E[6], i5F[6],
i60[6], i61[6], i62[6], i63[6], i64[6], i65[6], i66[6], i67[6],
i68[6], i69[6], i6A[6], i6B[6], i6C[6], i6D[6], i6E[6], i6F[6],
i70[6], i71[6], i72[6], i73[6], i74[6], i75[6], i76[6], i77[6],
i78[6], i79[6], i7A[6], i7B[6], i7C[6], i7D[6], i7E[6], i7F[6],
i80[6], i81[6], i82[6], i83[6], i84[6], i85[6], i86[6], i87[6],
i88[6], i89[6], i8A[6], i8B[6], i8C[6], i8D[6], i8E[6], i8F[6],
i90[6], i91[6], i92[6], i93[6], i94[6], i95[6], i96[6], i97[6],
i98[6], i99[6], i9A[6], i9B[6], i9C[6], i9D[6], i9E[6], i9F[6],
iA0[6], iA1[6], iA2[6], iA3[6], iA4[6], iA5[6], iA6[6], iA7[6],
iA8[6], iA9[6], iAA[6], iAB[6], iAC[6], iAD[6], iAE[6], iAF[6],
iB0[6], iB1[6], iB2[6], iB3[6], iB4[6], iB5[6], iB6[6], iB7[6],
iB8[6], iB9[6], iBA[6], iBB[6], iBC[6], iBD[6], iBE[6], iBF[6],
iC0[6], iC1[6], iC2[6], iC3[6], iC4[6], iC5[6], iC6[6], iC7[6],
iC8[6], iC9[6], iCA[6], iCB[6], iCC[6], iCD[6], iCE[6], iCF[6],
iD0[6], iD1[6], iD2[6], iD3[6], iD4[6], iD5[6], iD6[6], iD7[6],
iD8[6], iD9[6], iDA[6], iDB[6], iDC[6], iDD[6], iDE[6], iDF[6],
iE0[6], iE1[6], iE2[6], iE3[6], iE4[6], iE5[6], iE6[6], iE7[6],
iE8[6], iE9[6], iEA[6], iEB[6], iEC[6], iED[6], iEE[6], iEF[6],
iF0[6], iF1[6], iF2[6], iF3[6], iF4[6], iF5[6], iF6[6], iF7[6],
iF8[6], iF9[6], iFA[6], iFB[6], iFC[6], iFD[6], iFE[6], iFF[6]
}, S);


bitmux256 MX7(out[7], {
i00[7], i01[7], i02[7], i03[7], i04[7], i05[7], i06[7], i07[7],
i08[7], i09[7], i0A[7], i0B[7], i0C[7], i0D[7], i0E[7], i0F[7],
i10[7], i11[7], i12[7], i13[7], i14[7], i15[7], i16[7], i17[7],
i18[7], i19[7], i1A[7], i1B[7], i1C[7], i1D[7], i1E[7], i1F[7],
i20[7], i21[7], i22[7], i23[7], i24[7], i25[7], i26[7], i27[7],
i28[7], i29[7], i2A[7], i2B[7], i2C[7], i2D[7], i2E[7], i2F[7],
i30[7], i31[7], i32[7], i33[7], i34[7], i35[7], i36[7], i37[7],
i38[7], i39[7], i3A[7], i3B[7], i3C[7], i3D[7], i3E[7], i3F[7],
i40[7], i41[7], i42[7], i43[7], i44[7], i45[7], i46[7], i47[7],
i48[7], i49[7], i4A[7], i4B[7], i4C[7], i4D[7], i4E[7], i4F[7],
i50[7], i51[7], i52[7], i53[7], i54[7], i55[7], i56[7], i57[7],
i58[7], i59[7], i5A[7], i5B[7], i5C[7], i5D[7], i5E[7], i5F[7],
i60[7], i61[7], i62[7], i63[7], i64[7], i65[7], i66[7], i67[7],
i68[7], i69[7], i6A[7], i6B[7], i6C[7], i6D[7], i6E[7], i6F[7],
i70[7], i71[7], i72[7], i73[7], i74[7], i75[7], i76[7], i77[7],
i78[7], i79[7], i7A[7], i7B[7], i7C[7], i7D[7], i7E[7], i7F[7],
i80[7], i81[7], i82[7], i83[7], i84[7], i85[7], i86[7], i87[7],
i88[7], i89[7], i8A[7], i8B[7], i8C[7], i8D[7], i8E[7], i8F[7],
i90[7], i91[7], i92[7], i93[7], i94[7], i95[7], i96[7], i97[7],
i98[7], i99[7], i9A[7], i9B[7], i9C[7], i9D[7], i9E[7], i9F[7],
iA0[7], iA1[7], iA2[7], iA3[7], iA4[7], iA5[7], iA6[7], iA7[7],
iA8[7], iA9[7], iAA[7], iAB[7], iAC[7], iAD[7], iAE[7], iAF[7],
iB0[7], iB1[7], iB2[7], iB3[7], iB4[7], iB5[7], iB6[7], iB7[7],
iB8[7], iB9[7], iBA[7], iBB[7], iBC[7], iBD[7], iBE[7], iBF[7],
iC0[7], iC1[7], iC2[7], iC3[7], iC4[7], iC5[7], iC6[7], iC7[7],
iC8[7], iC9[7], iCA[7], iCB[7], iCC[7], iCD[7], iCE[7], iCF[7],
iD0[7], iD1[7], iD2[7], iD3[7], iD4[7], iD5[7], iD6[7], iD7[7],
iD8[7], iD9[7], iDA[7], iDB[7], iDC[7], iDD[7], iDE[7], iDF[7],
iE0[7], iE1[7], iE2[7], iE3[7], iE4[7], iE5[7], iE6[7], iE7[7],
iE8[7], iE9[7], iEA[7], iEB[7], iEC[7], iED[7], iEE[7], iEF[7],
iF0[7], iF1[7], iF2[7], iF3[7], iF4[7], iF5[7], iF6[7], iF7[7],
iF8[7], iF9[7], iFA[7], iFB[7], iFC[7], iFD[7], iFE[7], iFF[7]
}, S);


bitmux256 MX8(out[8], {
i00[8], i01[8], i02[8], i03[8], i04[8], i05[8], i06[8], i07[8],
i08[8], i09[8], i0A[8], i0B[8], i0C[8], i0D[8], i0E[8], i0F[8],
i10[8], i11[8], i12[8], i13[8], i14[8], i15[8], i16[8], i17[8],
i18[8], i19[8], i1A[8], i1B[8], i1C[8], i1D[8], i1E[8], i1F[8],
i20[8], i21[8], i22[8], i23[8], i24[8], i25[8], i26[8], i27[8],
i28[8], i29[8], i2A[8], i2B[8], i2C[8], i2D[8], i2E[8], i2F[8],
i30[8], i31[8], i32[8], i33[8], i34[8], i35[8], i36[8], i37[8],
i38[8], i39[8], i3A[8], i3B[8], i3C[8], i3D[8], i3E[8], i3F[8],
i40[8], i41[8], i42[8], i43[8], i44[8], i45[8], i46[8], i47[8],
i48[8], i49[8], i4A[8], i4B[8], i4C[8], i4D[8], i4E[8], i4F[8],
i50[8], i51[8], i52[8], i53[8], i54[8], i55[8], i56[8], i57[8],
i58[8], i59[8], i5A[8], i5B[8], i5C[8], i5D[8], i5E[8], i5F[8],
i60[8], i61[8], i62[8], i63[8], i64[8], i65[8], i66[8], i67[8],
i68[8], i69[8], i6A[8], i6B[8], i6C[8], i6D[8], i6E[8], i6F[8],
i70[8], i71[8], i72[8], i73[8], i74[8], i75[8], i76[8], i77[8],
i78[8], i79[8], i7A[8], i7B[8], i7C[8], i7D[8], i7E[8], i7F[8],
i80[8], i81[8], i82[8], i83[8], i84[8], i85[8], i86[8], i87[8],
i88[8], i89[8], i8A[8], i8B[8], i8C[8], i8D[8], i8E[8], i8F[8],
i90[8], i91[8], i92[8], i93[8], i94[8], i95[8], i96[8], i97[8],
i98[8], i99[8], i9A[8], i9B[8], i9C[8], i9D[8], i9E[8], i9F[8],
iA0[8], iA1[8], iA2[8], iA3[8], iA4[8], iA5[8], iA6[8], iA7[8],
iA8[8], iA9[8], iAA[8], iAB[8], iAC[8], iAD[8], iAE[8], iAF[8],
iB0[8], iB1[8], iB2[8], iB3[8], iB4[8], iB5[8], iB6[8], iB7[8],
iB8[8], iB9[8], iBA[8], iBB[8], iBC[8], iBD[8], iBE[8], iBF[8],
iC0[8], iC1[8], iC2[8], iC3[8], iC4[8], iC5[8], iC6[8], iC7[8],
iC8[8], iC9[8], iCA[8], iCB[8], iCC[8], iCD[8], iCE[8], iCF[8],
iD0[8], iD1[8], iD2[8], iD3[8], iD4[8], iD5[8], iD6[8], iD7[8],
iD8[8], iD9[8], iDA[8], iDB[8], iDC[8], iDD[8], iDE[8], iDF[8],
iE0[8], iE1[8], iE2[8], iE3[8], iE4[8], iE5[8], iE6[8], iE7[8],
iE8[8], iE9[8], iEA[8], iEB[8], iEC[8], iED[8], iEE[8], iEF[8],
iF0[8], iF1[8], iF2[8], iF3[8], iF4[8], iF5[8], iF6[8], iF7[8],
iF8[8], iF9[8], iFA[8], iFB[8], iFC[8], iFD[8], iFE[8], iFF[8]
}, S);


bitmux256 MX9(out[9], {
i00[9], i01[9], i02[9], i03[9], i04[9], i05[9], i06[9], i07[9],
i08[9], i09[9], i0A[9], i0B[9], i0C[9], i0D[9], i0E[9], i0F[9],
i10[9], i11[9], i12[9], i13[9], i14[9], i15[9], i16[9], i17[9],
i18[9], i19[9], i1A[9], i1B[9], i1C[9], i1D[9], i1E[9], i1F[9],
i20[9], i21[9], i22[9], i23[9], i24[9], i25[9], i26[9], i27[9],
i28[9], i29[9], i2A[9], i2B[9], i2C[9], i2D[9], i2E[9], i2F[9],
i30[9], i31[9], i32[9], i33[9], i34[9], i35[9], i36[9], i37[9],
i38[9], i39[9], i3A[9], i3B[9], i3C[9], i3D[9], i3E[9], i3F[9],
i40[9], i41[9], i42[9], i43[9], i44[9], i45[9], i46[9], i47[9],
i48[9], i49[9], i4A[9], i4B[9], i4C[9], i4D[9], i4E[9], i4F[9],
i50[9], i51[9], i52[9], i53[9], i54[9], i55[9], i56[9], i57[9],
i58[9], i59[9], i5A[9], i5B[9], i5C[9], i5D[9], i5E[9], i5F[9],
i60[9], i61[9], i62[9], i63[9], i64[9], i65[9], i66[9], i67[9],
i68[9], i69[9], i6A[9], i6B[9], i6C[9], i6D[9], i6E[9], i6F[9],
i70[9], i71[9], i72[9], i73[9], i74[9], i75[9], i76[9], i77[9],
i78[9], i79[9], i7A[9], i7B[9], i7C[9], i7D[9], i7E[9], i7F[9],
i80[9], i81[9], i82[9], i83[9], i84[9], i85[9], i86[9], i87[9],
i88[9], i89[9], i8A[9], i8B[9], i8C[9], i8D[9], i8E[9], i8F[9],
i90[9], i91[9], i92[9], i93[9], i94[9], i95[9], i96[9], i97[9],
i98[9], i99[9], i9A[9], i9B[9], i9C[9], i9D[9], i9E[9], i9F[9],
iA0[9], iA1[9], iA2[9], iA3[9], iA4[9], iA5[9], iA6[9], iA7[9],
iA8[9], iA9[9], iAA[9], iAB[9], iAC[9], iAD[9], iAE[9], iAF[9],
iB0[9], iB1[9], iB2[9], iB3[9], iB4[9], iB5[9], iB6[9], iB7[9],
iB8[9], iB9[9], iBA[9], iBB[9], iBC[9], iBD[9], iBE[9], iBF[9],
iC0[9], iC1[9], iC2[9], iC3[9], iC4[9], iC5[9], iC6[9], iC7[9],
iC8[9], iC9[9], iCA[9], iCB[9], iCC[9], iCD[9], iCE[9], iCF[9],
iD0[9], iD1[9], iD2[9], iD3[9], iD4[9], iD5[9], iD6[9], iD7[9],
iD8[9], iD9[9], iDA[9], iDB[9], iDC[9], iDD[9], iDE[9], iDF[9],
iE0[9], iE1[9], iE2[9], iE3[9], iE4[9], iE5[9], iE6[9], iE7[9],
iE8[9], iE9[9], iEA[9], iEB[9], iEC[9], iED[9], iEE[9], iEF[9],
iF0[9], iF1[9], iF2[9], iF3[9], iF4[9], iF5[9], iF6[9], iF7[9],
iF8[9], iF9[9], iFA[9], iFB[9], iFC[9], iFD[9], iFE[9], iFF[9]
}, S);


bitmux256 MX10(out[10], {
i00[10], i01[10], i02[10], i03[10], i04[10], i05[10], i06[10], i07[10],
i08[10], i09[10], i0A[10], i0B[10], i0C[10], i0D[10], i0E[10], i0F[10],
i10[10], i11[10], i12[10], i13[10], i14[10], i15[10], i16[10], i17[10],
i18[10], i19[10], i1A[10], i1B[10], i1C[10], i1D[10], i1E[10], i1F[10],
i20[10], i21[10], i22[10], i23[10], i24[10], i25[10], i26[10], i27[10],
i28[10], i29[10], i2A[10], i2B[10], i2C[10], i2D[10], i2E[10], i2F[10],
i30[10], i31[10], i32[10], i33[10], i34[10], i35[10], i36[10], i37[10],
i38[10], i39[10], i3A[10], i3B[10], i3C[10], i3D[10], i3E[10], i3F[10],
i40[10], i41[10], i42[10], i43[10], i44[10], i45[10], i46[10], i47[10],
i48[10], i49[10], i4A[10], i4B[10], i4C[10], i4D[10], i4E[10], i4F[10],
i50[10], i51[10], i52[10], i53[10], i54[10], i55[10], i56[10], i57[10],
i58[10], i59[10], i5A[10], i5B[10], i5C[10], i5D[10], i5E[10], i5F[10],
i60[10], i61[10], i62[10], i63[10], i64[10], i65[10], i66[10], i67[10],
i68[10], i69[10], i6A[10], i6B[10], i6C[10], i6D[10], i6E[10], i6F[10],
i70[10], i71[10], i72[10], i73[10], i74[10], i75[10], i76[10], i77[10],
i78[10], i79[10], i7A[10], i7B[10], i7C[10], i7D[10], i7E[10], i7F[10],
i80[10], i81[10], i82[10], i83[10], i84[10], i85[10], i86[10], i87[10],
i88[10], i89[10], i8A[10], i8B[10], i8C[10], i8D[10], i8E[10], i8F[10],
i90[10], i91[10], i92[10], i93[10], i94[10], i95[10], i96[10], i97[10],
i98[10], i99[10], i9A[10], i9B[10], i9C[10], i9D[10], i9E[10], i9F[10],
iA0[10], iA1[10], iA2[10], iA3[10], iA4[10], iA5[10], iA6[10], iA7[10],
iA8[10], iA9[10], iAA[10], iAB[10], iAC[10], iAD[10], iAE[10], iAF[10],
iB0[10], iB1[10], iB2[10], iB3[10], iB4[10], iB5[10], iB6[10], iB7[10],
iB8[10], iB9[10], iBA[10], iBB[10], iBC[10], iBD[10], iBE[10], iBF[10],
iC0[10], iC1[10], iC2[10], iC3[10], iC4[10], iC5[10], iC6[10], iC7[10],
iC8[10], iC9[10], iCA[10], iCB[10], iCC[10], iCD[10], iCE[10], iCF[10],
iD0[10], iD1[10], iD2[10], iD3[10], iD4[10], iD5[10], iD6[10], iD7[10],
iD8[10], iD9[10], iDA[10], iDB[10], iDC[10], iDD[10], iDE[10], iDF[10],
iE0[10], iE1[10], iE2[10], iE3[10], iE4[10], iE5[10], iE6[10], iE7[10],
iE8[10], iE9[10], iEA[10], iEB[10], iEC[10], iED[10], iEE[10], iEF[10],
iF0[10], iF1[10], iF2[10], iF3[10], iF4[10], iF5[10], iF6[10], iF7[10],
iF8[10], iF9[10], iFA[10], iFB[10], iFC[10], iFD[10], iFE[10], iFF[10]
}, S);


bitmux256 MX11(out[11], {
i00[11], i01[11], i02[11], i03[11], i04[11], i05[11], i06[11], i07[11],
i08[11], i09[11], i0A[11], i0B[11], i0C[11], i0D[11], i0E[11], i0F[11],
i10[11], i11[11], i12[11], i13[11], i14[11], i15[11], i16[11], i17[11],
i18[11], i19[11], i1A[11], i1B[11], i1C[11], i1D[11], i1E[11], i1F[11],
i20[11], i21[11], i22[11], i23[11], i24[11], i25[11], i26[11], i27[11],
i28[11], i29[11], i2A[11], i2B[11], i2C[11], i2D[11], i2E[11], i2F[11],
i30[11], i31[11], i32[11], i33[11], i34[11], i35[11], i36[11], i37[11],
i38[11], i39[11], i3A[11], i3B[11], i3C[11], i3D[11], i3E[11], i3F[11],
i40[11], i41[11], i42[11], i43[11], i44[11], i45[11], i46[11], i47[11],
i48[11], i49[11], i4A[11], i4B[11], i4C[11], i4D[11], i4E[11], i4F[11],
i50[11], i51[11], i52[11], i53[11], i54[11], i55[11], i56[11], i57[11],
i58[11], i59[11], i5A[11], i5B[11], i5C[11], i5D[11], i5E[11], i5F[11],
i60[11], i61[11], i62[11], i63[11], i64[11], i65[11], i66[11], i67[11],
i68[11], i69[11], i6A[11], i6B[11], i6C[11], i6D[11], i6E[11], i6F[11],
i70[11], i71[11], i72[11], i73[11], i74[11], i75[11], i76[11], i77[11],
i78[11], i79[11], i7A[11], i7B[11], i7C[11], i7D[11], i7E[11], i7F[11],
i80[11], i81[11], i82[11], i83[11], i84[11], i85[11], i86[11], i87[11],
i88[11], i89[11], i8A[11], i8B[11], i8C[11], i8D[11], i8E[11], i8F[11],
i90[11], i91[11], i92[11], i93[11], i94[11], i95[11], i96[11], i97[11],
i98[11], i99[11], i9A[11], i9B[11], i9C[11], i9D[11], i9E[11], i9F[11],
iA0[11], iA1[11], iA2[11], iA3[11], iA4[11], iA5[11], iA6[11], iA7[11],
iA8[11], iA9[11], iAA[11], iAB[11], iAC[11], iAD[11], iAE[11], iAF[11],
iB0[11], iB1[11], iB2[11], iB3[11], iB4[11], iB5[11], iB6[11], iB7[11],
iB8[11], iB9[11], iBA[11], iBB[11], iBC[11], iBD[11], iBE[11], iBF[11],
iC0[11], iC1[11], iC2[11], iC3[11], iC4[11], iC5[11], iC6[11], iC7[11],
iC8[11], iC9[11], iCA[11], iCB[11], iCC[11], iCD[11], iCE[11], iCF[11],
iD0[11], iD1[11], iD2[11], iD3[11], iD4[11], iD5[11], iD6[11], iD7[11],
iD8[11], iD9[11], iDA[11], iDB[11], iDC[11], iDD[11], iDE[11], iDF[11],
iE0[11], iE1[11], iE2[11], iE3[11], iE4[11], iE5[11], iE6[11], iE7[11],
iE8[11], iE9[11], iEA[11], iEB[11], iEC[11], iED[11], iEE[11], iEF[11],
iF0[11], iF1[11], iF2[11], iF3[11], iF4[11], iF5[11], iF6[11], iF7[11],
iF8[11], iF9[11], iFA[11], iFB[11], iFC[11], iFD[11], iFE[11], iFF[11]
}, S);


bitmux256 MX12(out[12], {
i00[12], i01[12], i02[12], i03[12], i04[12], i05[12], i06[12], i07[12],
i08[12], i09[12], i0A[12], i0B[12], i0C[12], i0D[12], i0E[12], i0F[12],
i10[12], i11[12], i12[12], i13[12], i14[12], i15[12], i16[12], i17[12],
i18[12], i19[12], i1A[12], i1B[12], i1C[12], i1D[12], i1E[12], i1F[12],
i20[12], i21[12], i22[12], i23[12], i24[12], i25[12], i26[12], i27[12],
i28[12], i29[12], i2A[12], i2B[12], i2C[12], i2D[12], i2E[12], i2F[12],
i30[12], i31[12], i32[12], i33[12], i34[12], i35[12], i36[12], i37[12],
i38[12], i39[12], i3A[12], i3B[12], i3C[12], i3D[12], i3E[12], i3F[12],
i40[12], i41[12], i42[12], i43[12], i44[12], i45[12], i46[12], i47[12],
i48[12], i49[12], i4A[12], i4B[12], i4C[12], i4D[12], i4E[12], i4F[12],
i50[12], i51[12], i52[12], i53[12], i54[12], i55[12], i56[12], i57[12],
i58[12], i59[12], i5A[12], i5B[12], i5C[12], i5D[12], i5E[12], i5F[12],
i60[12], i61[12], i62[12], i63[12], i64[12], i65[12], i66[12], i67[12],
i68[12], i69[12], i6A[12], i6B[12], i6C[12], i6D[12], i6E[12], i6F[12],
i70[12], i71[12], i72[12], i73[12], i74[12], i75[12], i76[12], i77[12],
i78[12], i79[12], i7A[12], i7B[12], i7C[12], i7D[12], i7E[12], i7F[12],
i80[12], i81[12], i82[12], i83[12], i84[12], i85[12], i86[12], i87[12],
i88[12], i89[12], i8A[12], i8B[12], i8C[12], i8D[12], i8E[12], i8F[12],
i90[12], i91[12], i92[12], i93[12], i94[12], i95[12], i96[12], i97[12],
i98[12], i99[12], i9A[12], i9B[12], i9C[12], i9D[12], i9E[12], i9F[12],
iA0[12], iA1[12], iA2[12], iA3[12], iA4[12], iA5[12], iA6[12], iA7[12],
iA8[12], iA9[12], iAA[12], iAB[12], iAC[12], iAD[12], iAE[12], iAF[12],
iB0[12], iB1[12], iB2[12], iB3[12], iB4[12], iB5[12], iB6[12], iB7[12],
iB8[12], iB9[12], iBA[12], iBB[12], iBC[12], iBD[12], iBE[12], iBF[12],
iC0[12], iC1[12], iC2[12], iC3[12], iC4[12], iC5[12], iC6[12], iC7[12],
iC8[12], iC9[12], iCA[12], iCB[12], iCC[12], iCD[12], iCE[12], iCF[12],
iD0[12], iD1[12], iD2[12], iD3[12], iD4[12], iD5[12], iD6[12], iD7[12],
iD8[12], iD9[12], iDA[12], iDB[12], iDC[12], iDD[12], iDE[12], iDF[12],
iE0[12], iE1[12], iE2[12], iE3[12], iE4[12], iE5[12], iE6[12], iE7[12],
iE8[12], iE9[12], iEA[12], iEB[12], iEC[12], iED[12], iEE[12], iEF[12],
iF0[12], iF1[12], iF2[12], iF3[12], iF4[12], iF5[12], iF6[12], iF7[12],
iF8[12], iF9[12], iFA[12], iFB[12], iFC[12], iFD[12], iFE[12], iFF[12]
}, S);


bitmux256 MX13(out[13], {
i00[13], i01[13], i02[13], i03[13], i04[13], i05[13], i06[13], i07[13],
i08[13], i09[13], i0A[13], i0B[13], i0C[13], i0D[13], i0E[13], i0F[13],
i10[13], i11[13], i12[13], i13[13], i14[13], i15[13], i16[13], i17[13],
i18[13], i19[13], i1A[13], i1B[13], i1C[13], i1D[13], i1E[13], i1F[13],
i20[13], i21[13], i22[13], i23[13], i24[13], i25[13], i26[13], i27[13],
i28[13], i29[13], i2A[13], i2B[13], i2C[13], i2D[13], i2E[13], i2F[13],
i30[13], i31[13], i32[13], i33[13], i34[13], i35[13], i36[13], i37[13],
i38[13], i39[13], i3A[13], i3B[13], i3C[13], i3D[13], i3E[13], i3F[13],
i40[13], i41[13], i42[13], i43[13], i44[13], i45[13], i46[13], i47[13],
i48[13], i49[13], i4A[13], i4B[13], i4C[13], i4D[13], i4E[13], i4F[13],
i50[13], i51[13], i52[13], i53[13], i54[13], i55[13], i56[13], i57[13],
i58[13], i59[13], i5A[13], i5B[13], i5C[13], i5D[13], i5E[13], i5F[13],
i60[13], i61[13], i62[13], i63[13], i64[13], i65[13], i66[13], i67[13],
i68[13], i69[13], i6A[13], i6B[13], i6C[13], i6D[13], i6E[13], i6F[13],
i70[13], i71[13], i72[13], i73[13], i74[13], i75[13], i76[13], i77[13],
i78[13], i79[13], i7A[13], i7B[13], i7C[13], i7D[13], i7E[13], i7F[13],
i80[13], i81[13], i82[13], i83[13], i84[13], i85[13], i86[13], i87[13],
i88[13], i89[13], i8A[13], i8B[13], i8C[13], i8D[13], i8E[13], i8F[13],
i90[13], i91[13], i92[13], i93[13], i94[13], i95[13], i96[13], i97[13],
i98[13], i99[13], i9A[13], i9B[13], i9C[13], i9D[13], i9E[13], i9F[13],
iA0[13], iA1[13], iA2[13], iA3[13], iA4[13], iA5[13], iA6[13], iA7[13],
iA8[13], iA9[13], iAA[13], iAB[13], iAC[13], iAD[13], iAE[13], iAF[13],
iB0[13], iB1[13], iB2[13], iB3[13], iB4[13], iB5[13], iB6[13], iB7[13],
iB8[13], iB9[13], iBA[13], iBB[13], iBC[13], iBD[13], iBE[13], iBF[13],
iC0[13], iC1[13], iC2[13], iC3[13], iC4[13], iC5[13], iC6[13], iC7[13],
iC8[13], iC9[13], iCA[13], iCB[13], iCC[13], iCD[13], iCE[13], iCF[13],
iD0[13], iD1[13], iD2[13], iD3[13], iD4[13], iD5[13], iD6[13], iD7[13],
iD8[13], iD9[13], iDA[13], iDB[13], iDC[13], iDD[13], iDE[13], iDF[13],
iE0[13], iE1[13], iE2[13], iE3[13], iE4[13], iE5[13], iE6[13], iE7[13],
iE8[13], iE9[13], iEA[13], iEB[13], iEC[13], iED[13], iEE[13], iEF[13],
iF0[13], iF1[13], iF2[13], iF3[13], iF4[13], iF5[13], iF6[13], iF7[13],
iF8[13], iF9[13], iFA[13], iFB[13], iFC[13], iFD[13], iFE[13], iFF[13]
}, S);


bitmux256 MX14(out[14], {
i00[14], i01[14], i02[14], i03[14], i04[14], i05[14], i06[14], i07[14],
i08[14], i09[14], i0A[14], i0B[14], i0C[14], i0D[14], i0E[14], i0F[14],
i10[14], i11[14], i12[14], i13[14], i14[14], i15[14], i16[14], i17[14],
i18[14], i19[14], i1A[14], i1B[14], i1C[14], i1D[14], i1E[14], i1F[14],
i20[14], i21[14], i22[14], i23[14], i24[14], i25[14], i26[14], i27[14],
i28[14], i29[14], i2A[14], i2B[14], i2C[14], i2D[14], i2E[14], i2F[14],
i30[14], i31[14], i32[14], i33[14], i34[14], i35[14], i36[14], i37[14],
i38[14], i39[14], i3A[14], i3B[14], i3C[14], i3D[14], i3E[14], i3F[14],
i40[14], i41[14], i42[14], i43[14], i44[14], i45[14], i46[14], i47[14],
i48[14], i49[14], i4A[14], i4B[14], i4C[14], i4D[14], i4E[14], i4F[14],
i50[14], i51[14], i52[14], i53[14], i54[14], i55[14], i56[14], i57[14],
i58[14], i59[14], i5A[14], i5B[14], i5C[14], i5D[14], i5E[14], i5F[14],
i60[14], i61[14], i62[14], i63[14], i64[14], i65[14], i66[14], i67[14],
i68[14], i69[14], i6A[14], i6B[14], i6C[14], i6D[14], i6E[14], i6F[14],
i70[14], i71[14], i72[14], i73[14], i74[14], i75[14], i76[14], i77[14],
i78[14], i79[14], i7A[14], i7B[14], i7C[14], i7D[14], i7E[14], i7F[14],
i80[14], i81[14], i82[14], i83[14], i84[14], i85[14], i86[14], i87[14],
i88[14], i89[14], i8A[14], i8B[14], i8C[14], i8D[14], i8E[14], i8F[14],
i90[14], i91[14], i92[14], i93[14], i94[14], i95[14], i96[14], i97[14],
i98[14], i99[14], i9A[14], i9B[14], i9C[14], i9D[14], i9E[14], i9F[14],
iA0[14], iA1[14], iA2[14], iA3[14], iA4[14], iA5[14], iA6[14], iA7[14],
iA8[14], iA9[14], iAA[14], iAB[14], iAC[14], iAD[14], iAE[14], iAF[14],
iB0[14], iB1[14], iB2[14], iB3[14], iB4[14], iB5[14], iB6[14], iB7[14],
iB8[14], iB9[14], iBA[14], iBB[14], iBC[14], iBD[14], iBE[14], iBF[14],
iC0[14], iC1[14], iC2[14], iC3[14], iC4[14], iC5[14], iC6[14], iC7[14],
iC8[14], iC9[14], iCA[14], iCB[14], iCC[14], iCD[14], iCE[14], iCF[14],
iD0[14], iD1[14], iD2[14], iD3[14], iD4[14], iD5[14], iD6[14], iD7[14],
iD8[14], iD9[14], iDA[14], iDB[14], iDC[14], iDD[14], iDE[14], iDF[14],
iE0[14], iE1[14], iE2[14], iE3[14], iE4[14], iE5[14], iE6[14], iE7[14],
iE8[14], iE9[14], iEA[14], iEB[14], iEC[14], iED[14], iEE[14], iEF[14],
iF0[14], iF1[14], iF2[14], iF3[14], iF4[14], iF5[14], iF6[14], iF7[14],
iF8[14], iF9[14], iFA[14], iFB[14], iFC[14], iFD[14], iFE[14], iFF[14]
}, S);


bitmux256 MX15(out[15], {
i00[15], i01[15], i02[15], i03[15], i04[15], i05[15], i06[15], i07[15],
i08[15], i09[15], i0A[15], i0B[15], i0C[15], i0D[15], i0E[15], i0F[15],
i10[15], i11[15], i12[15], i13[15], i14[15], i15[15], i16[15], i17[15],
i18[15], i19[15], i1A[15], i1B[15], i1C[15], i1D[15], i1E[15], i1F[15],
i20[15], i21[15], i22[15], i23[15], i24[15], i25[15], i26[15], i27[15],
i28[15], i29[15], i2A[15], i2B[15], i2C[15], i2D[15], i2E[15], i2F[15],
i30[15], i31[15], i32[15], i33[15], i34[15], i35[15], i36[15], i37[15],
i38[15], i39[15], i3A[15], i3B[15], i3C[15], i3D[15], i3E[15], i3F[15],
i40[15], i41[15], i42[15], i43[15], i44[15], i45[15], i46[15], i47[15],
i48[15], i49[15], i4A[15], i4B[15], i4C[15], i4D[15], i4E[15], i4F[15],
i50[15], i51[15], i52[15], i53[15], i54[15], i55[15], i56[15], i57[15],
i58[15], i59[15], i5A[15], i5B[15], i5C[15], i5D[15], i5E[15], i5F[15],
i60[15], i61[15], i62[15], i63[15], i64[15], i65[15], i66[15], i67[15],
i68[15], i69[15], i6A[15], i6B[15], i6C[15], i6D[15], i6E[15], i6F[15],
i70[15], i71[15], i72[15], i73[15], i74[15], i75[15], i76[15], i77[15],
i78[15], i79[15], i7A[15], i7B[15], i7C[15], i7D[15], i7E[15], i7F[15],
i80[15], i81[15], i82[15], i83[15], i84[15], i85[15], i86[15], i87[15],
i88[15], i89[15], i8A[15], i8B[15], i8C[15], i8D[15], i8E[15], i8F[15],
i90[15], i91[15], i92[15], i93[15], i94[15], i95[15], i96[15], i97[15],
i98[15], i99[15], i9A[15], i9B[15], i9C[15], i9D[15], i9E[15], i9F[15],
iA0[15], iA1[15], iA2[15], iA3[15], iA4[15], iA5[15], iA6[15], iA7[15],
iA8[15], iA9[15], iAA[15], iAB[15], iAC[15], iAD[15], iAE[15], iAF[15],
iB0[15], iB1[15], iB2[15], iB3[15], iB4[15], iB5[15], iB6[15], iB7[15],
iB8[15], iB9[15], iBA[15], iBB[15], iBC[15], iBD[15], iBE[15], iBF[15],
iC0[15], iC1[15], iC2[15], iC3[15], iC4[15], iC5[15], iC6[15], iC7[15],
iC8[15], iC9[15], iCA[15], iCB[15], iCC[15], iCD[15], iCE[15], iCF[15],
iD0[15], iD1[15], iD2[15], iD3[15], iD4[15], iD5[15], iD6[15], iD7[15],
iD8[15], iD9[15], iDA[15], iDB[15], iDC[15], iDD[15], iDE[15], iDF[15],
iE0[15], iE1[15], iE2[15], iE3[15], iE4[15], iE5[15], iE6[15], iE7[15],
iE8[15], iE9[15], iEA[15], iEB[15], iEC[15], iED[15], iEE[15], iEF[15],
iF0[15], iF1[15], iF2[15], iF3[15], iF4[15], iF5[15], iF6[15], iF7[15],
iF8[15], iF9[15], iFA[15], iFB[15], iFC[15], iFD[15], iFE[15], iFF[15]
}, S);


bitmux256 MX16(out[16], {
i00[16], i01[16], i02[16], i03[16], i04[16], i05[16], i06[16], i07[16],
i08[16], i09[16], i0A[16], i0B[16], i0C[16], i0D[16], i0E[16], i0F[16],
i10[16], i11[16], i12[16], i13[16], i14[16], i15[16], i16[16], i17[16],
i18[16], i19[16], i1A[16], i1B[16], i1C[16], i1D[16], i1E[16], i1F[16],
i20[16], i21[16], i22[16], i23[16], i24[16], i25[16], i26[16], i27[16],
i28[16], i29[16], i2A[16], i2B[16], i2C[16], i2D[16], i2E[16], i2F[16],
i30[16], i31[16], i32[16], i33[16], i34[16], i35[16], i36[16], i37[16],
i38[16], i39[16], i3A[16], i3B[16], i3C[16], i3D[16], i3E[16], i3F[16],
i40[16], i41[16], i42[16], i43[16], i44[16], i45[16], i46[16], i47[16],
i48[16], i49[16], i4A[16], i4B[16], i4C[16], i4D[16], i4E[16], i4F[16],
i50[16], i51[16], i52[16], i53[16], i54[16], i55[16], i56[16], i57[16],
i58[16], i59[16], i5A[16], i5B[16], i5C[16], i5D[16], i5E[16], i5F[16],
i60[16], i61[16], i62[16], i63[16], i64[16], i65[16], i66[16], i67[16],
i68[16], i69[16], i6A[16], i6B[16], i6C[16], i6D[16], i6E[16], i6F[16],
i70[16], i71[16], i72[16], i73[16], i74[16], i75[16], i76[16], i77[16],
i78[16], i79[16], i7A[16], i7B[16], i7C[16], i7D[16], i7E[16], i7F[16],
i80[16], i81[16], i82[16], i83[16], i84[16], i85[16], i86[16], i87[16],
i88[16], i89[16], i8A[16], i8B[16], i8C[16], i8D[16], i8E[16], i8F[16],
i90[16], i91[16], i92[16], i93[16], i94[16], i95[16], i96[16], i97[16],
i98[16], i99[16], i9A[16], i9B[16], i9C[16], i9D[16], i9E[16], i9F[16],
iA0[16], iA1[16], iA2[16], iA3[16], iA4[16], iA5[16], iA6[16], iA7[16],
iA8[16], iA9[16], iAA[16], iAB[16], iAC[16], iAD[16], iAE[16], iAF[16],
iB0[16], iB1[16], iB2[16], iB3[16], iB4[16], iB5[16], iB6[16], iB7[16],
iB8[16], iB9[16], iBA[16], iBB[16], iBC[16], iBD[16], iBE[16], iBF[16],
iC0[16], iC1[16], iC2[16], iC3[16], iC4[16], iC5[16], iC6[16], iC7[16],
iC8[16], iC9[16], iCA[16], iCB[16], iCC[16], iCD[16], iCE[16], iCF[16],
iD0[16], iD1[16], iD2[16], iD3[16], iD4[16], iD5[16], iD6[16], iD7[16],
iD8[16], iD9[16], iDA[16], iDB[16], iDC[16], iDD[16], iDE[16], iDF[16],
iE0[16], iE1[16], iE2[16], iE3[16], iE4[16], iE5[16], iE6[16], iE7[16],
iE8[16], iE9[16], iEA[16], iEB[16], iEC[16], iED[16], iEE[16], iEF[16],
iF0[16], iF1[16], iF2[16], iF3[16], iF4[16], iF5[16], iF6[16], iF7[16],
iF8[16], iF9[16], iFA[16], iFB[16], iFC[16], iFD[16], iFE[16], iFF[16]
}, S);


bitmux256 MX17(out[17], {
i00[17], i01[17], i02[17], i03[17], i04[17], i05[17], i06[17], i07[17],
i08[17], i09[17], i0A[17], i0B[17], i0C[17], i0D[17], i0E[17], i0F[17],
i10[17], i11[17], i12[17], i13[17], i14[17], i15[17], i16[17], i17[17],
i18[17], i19[17], i1A[17], i1B[17], i1C[17], i1D[17], i1E[17], i1F[17],
i20[17], i21[17], i22[17], i23[17], i24[17], i25[17], i26[17], i27[17],
i28[17], i29[17], i2A[17], i2B[17], i2C[17], i2D[17], i2E[17], i2F[17],
i30[17], i31[17], i32[17], i33[17], i34[17], i35[17], i36[17], i37[17],
i38[17], i39[17], i3A[17], i3B[17], i3C[17], i3D[17], i3E[17], i3F[17],
i40[17], i41[17], i42[17], i43[17], i44[17], i45[17], i46[17], i47[17],
i48[17], i49[17], i4A[17], i4B[17], i4C[17], i4D[17], i4E[17], i4F[17],
i50[17], i51[17], i52[17], i53[17], i54[17], i55[17], i56[17], i57[17],
i58[17], i59[17], i5A[17], i5B[17], i5C[17], i5D[17], i5E[17], i5F[17],
i60[17], i61[17], i62[17], i63[17], i64[17], i65[17], i66[17], i67[17],
i68[17], i69[17], i6A[17], i6B[17], i6C[17], i6D[17], i6E[17], i6F[17],
i70[17], i71[17], i72[17], i73[17], i74[17], i75[17], i76[17], i77[17],
i78[17], i79[17], i7A[17], i7B[17], i7C[17], i7D[17], i7E[17], i7F[17],
i80[17], i81[17], i82[17], i83[17], i84[17], i85[17], i86[17], i87[17],
i88[17], i89[17], i8A[17], i8B[17], i8C[17], i8D[17], i8E[17], i8F[17],
i90[17], i91[17], i92[17], i93[17], i94[17], i95[17], i96[17], i97[17],
i98[17], i99[17], i9A[17], i9B[17], i9C[17], i9D[17], i9E[17], i9F[17],
iA0[17], iA1[17], iA2[17], iA3[17], iA4[17], iA5[17], iA6[17], iA7[17],
iA8[17], iA9[17], iAA[17], iAB[17], iAC[17], iAD[17], iAE[17], iAF[17],
iB0[17], iB1[17], iB2[17], iB3[17], iB4[17], iB5[17], iB6[17], iB7[17],
iB8[17], iB9[17], iBA[17], iBB[17], iBC[17], iBD[17], iBE[17], iBF[17],
iC0[17], iC1[17], iC2[17], iC3[17], iC4[17], iC5[17], iC6[17], iC7[17],
iC8[17], iC9[17], iCA[17], iCB[17], iCC[17], iCD[17], iCE[17], iCF[17],
iD0[17], iD1[17], iD2[17], iD3[17], iD4[17], iD5[17], iD6[17], iD7[17],
iD8[17], iD9[17], iDA[17], iDB[17], iDC[17], iDD[17], iDE[17], iDF[17],
iE0[17], iE1[17], iE2[17], iE3[17], iE4[17], iE5[17], iE6[17], iE7[17],
iE8[17], iE9[17], iEA[17], iEB[17], iEC[17], iED[17], iEE[17], iEF[17],
iF0[17], iF1[17], iF2[17], iF3[17], iF4[17], iF5[17], iF6[17], iF7[17],
iF8[17], iF9[17], iFA[17], iFB[17], iFC[17], iFD[17], iFE[17], iFF[17]
}, S);


bitmux256 MX18(out[18], {
i00[18], i01[18], i02[18], i03[18], i04[18], i05[18], i06[18], i07[18],
i08[18], i09[18], i0A[18], i0B[18], i0C[18], i0D[18], i0E[18], i0F[18],
i10[18], i11[18], i12[18], i13[18], i14[18], i15[18], i16[18], i17[18],
i18[18], i19[18], i1A[18], i1B[18], i1C[18], i1D[18], i1E[18], i1F[18],
i20[18], i21[18], i22[18], i23[18], i24[18], i25[18], i26[18], i27[18],
i28[18], i29[18], i2A[18], i2B[18], i2C[18], i2D[18], i2E[18], i2F[18],
i30[18], i31[18], i32[18], i33[18], i34[18], i35[18], i36[18], i37[18],
i38[18], i39[18], i3A[18], i3B[18], i3C[18], i3D[18], i3E[18], i3F[18],
i40[18], i41[18], i42[18], i43[18], i44[18], i45[18], i46[18], i47[18],
i48[18], i49[18], i4A[18], i4B[18], i4C[18], i4D[18], i4E[18], i4F[18],
i50[18], i51[18], i52[18], i53[18], i54[18], i55[18], i56[18], i57[18],
i58[18], i59[18], i5A[18], i5B[18], i5C[18], i5D[18], i5E[18], i5F[18],
i60[18], i61[18], i62[18], i63[18], i64[18], i65[18], i66[18], i67[18],
i68[18], i69[18], i6A[18], i6B[18], i6C[18], i6D[18], i6E[18], i6F[18],
i70[18], i71[18], i72[18], i73[18], i74[18], i75[18], i76[18], i77[18],
i78[18], i79[18], i7A[18], i7B[18], i7C[18], i7D[18], i7E[18], i7F[18],
i80[18], i81[18], i82[18], i83[18], i84[18], i85[18], i86[18], i87[18],
i88[18], i89[18], i8A[18], i8B[18], i8C[18], i8D[18], i8E[18], i8F[18],
i90[18], i91[18], i92[18], i93[18], i94[18], i95[18], i96[18], i97[18],
i98[18], i99[18], i9A[18], i9B[18], i9C[18], i9D[18], i9E[18], i9F[18],
iA0[18], iA1[18], iA2[18], iA3[18], iA4[18], iA5[18], iA6[18], iA7[18],
iA8[18], iA9[18], iAA[18], iAB[18], iAC[18], iAD[18], iAE[18], iAF[18],
iB0[18], iB1[18], iB2[18], iB3[18], iB4[18], iB5[18], iB6[18], iB7[18],
iB8[18], iB9[18], iBA[18], iBB[18], iBC[18], iBD[18], iBE[18], iBF[18],
iC0[18], iC1[18], iC2[18], iC3[18], iC4[18], iC5[18], iC6[18], iC7[18],
iC8[18], iC9[18], iCA[18], iCB[18], iCC[18], iCD[18], iCE[18], iCF[18],
iD0[18], iD1[18], iD2[18], iD3[18], iD4[18], iD5[18], iD6[18], iD7[18],
iD8[18], iD9[18], iDA[18], iDB[18], iDC[18], iDD[18], iDE[18], iDF[18],
iE0[18], iE1[18], iE2[18], iE3[18], iE4[18], iE5[18], iE6[18], iE7[18],
iE8[18], iE9[18], iEA[18], iEB[18], iEC[18], iED[18], iEE[18], iEF[18],
iF0[18], iF1[18], iF2[18], iF3[18], iF4[18], iF5[18], iF6[18], iF7[18],
iF8[18], iF9[18], iFA[18], iFB[18], iFC[18], iFD[18], iFE[18], iFF[18]
}, S);


bitmux256 MX19(out[19], {
i00[19], i01[19], i02[19], i03[19], i04[19], i05[19], i06[19], i07[19],
i08[19], i09[19], i0A[19], i0B[19], i0C[19], i0D[19], i0E[19], i0F[19],
i10[19], i11[19], i12[19], i13[19], i14[19], i15[19], i16[19], i17[19],
i18[19], i19[19], i1A[19], i1B[19], i1C[19], i1D[19], i1E[19], i1F[19],
i20[19], i21[19], i22[19], i23[19], i24[19], i25[19], i26[19], i27[19],
i28[19], i29[19], i2A[19], i2B[19], i2C[19], i2D[19], i2E[19], i2F[19],
i30[19], i31[19], i32[19], i33[19], i34[19], i35[19], i36[19], i37[19],
i38[19], i39[19], i3A[19], i3B[19], i3C[19], i3D[19], i3E[19], i3F[19],
i40[19], i41[19], i42[19], i43[19], i44[19], i45[19], i46[19], i47[19],
i48[19], i49[19], i4A[19], i4B[19], i4C[19], i4D[19], i4E[19], i4F[19],
i50[19], i51[19], i52[19], i53[19], i54[19], i55[19], i56[19], i57[19],
i58[19], i59[19], i5A[19], i5B[19], i5C[19], i5D[19], i5E[19], i5F[19],
i60[19], i61[19], i62[19], i63[19], i64[19], i65[19], i66[19], i67[19],
i68[19], i69[19], i6A[19], i6B[19], i6C[19], i6D[19], i6E[19], i6F[19],
i70[19], i71[19], i72[19], i73[19], i74[19], i75[19], i76[19], i77[19],
i78[19], i79[19], i7A[19], i7B[19], i7C[19], i7D[19], i7E[19], i7F[19],
i80[19], i81[19], i82[19], i83[19], i84[19], i85[19], i86[19], i87[19],
i88[19], i89[19], i8A[19], i8B[19], i8C[19], i8D[19], i8E[19], i8F[19],
i90[19], i91[19], i92[19], i93[19], i94[19], i95[19], i96[19], i97[19],
i98[19], i99[19], i9A[19], i9B[19], i9C[19], i9D[19], i9E[19], i9F[19],
iA0[19], iA1[19], iA2[19], iA3[19], iA4[19], iA5[19], iA6[19], iA7[19],
iA8[19], iA9[19], iAA[19], iAB[19], iAC[19], iAD[19], iAE[19], iAF[19],
iB0[19], iB1[19], iB2[19], iB3[19], iB4[19], iB5[19], iB6[19], iB7[19],
iB8[19], iB9[19], iBA[19], iBB[19], iBC[19], iBD[19], iBE[19], iBF[19],
iC0[19], iC1[19], iC2[19], iC3[19], iC4[19], iC5[19], iC6[19], iC7[19],
iC8[19], iC9[19], iCA[19], iCB[19], iCC[19], iCD[19], iCE[19], iCF[19],
iD0[19], iD1[19], iD2[19], iD3[19], iD4[19], iD5[19], iD6[19], iD7[19],
iD8[19], iD9[19], iDA[19], iDB[19], iDC[19], iDD[19], iDE[19], iDF[19],
iE0[19], iE1[19], iE2[19], iE3[19], iE4[19], iE5[19], iE6[19], iE7[19],
iE8[19], iE9[19], iEA[19], iEB[19], iEC[19], iED[19], iEE[19], iEF[19],
iF0[19], iF1[19], iF2[19], iF3[19], iF4[19], iF5[19], iF6[19], iF7[19],
iF8[19], iF9[19], iFA[19], iFB[19], iFC[19], iFD[19], iFE[19], iFF[19]
}, S);


bitmux256 MX20(out[20], {
i00[20], i01[20], i02[20], i03[20], i04[20], i05[20], i06[20], i07[20],
i08[20], i09[20], i0A[20], i0B[20], i0C[20], i0D[20], i0E[20], i0F[20],
i10[20], i11[20], i12[20], i13[20], i14[20], i15[20], i16[20], i17[20],
i18[20], i19[20], i1A[20], i1B[20], i1C[20], i1D[20], i1E[20], i1F[20],
i20[20], i21[20], i22[20], i23[20], i24[20], i25[20], i26[20], i27[20],
i28[20], i29[20], i2A[20], i2B[20], i2C[20], i2D[20], i2E[20], i2F[20],
i30[20], i31[20], i32[20], i33[20], i34[20], i35[20], i36[20], i37[20],
i38[20], i39[20], i3A[20], i3B[20], i3C[20], i3D[20], i3E[20], i3F[20],
i40[20], i41[20], i42[20], i43[20], i44[20], i45[20], i46[20], i47[20],
i48[20], i49[20], i4A[20], i4B[20], i4C[20], i4D[20], i4E[20], i4F[20],
i50[20], i51[20], i52[20], i53[20], i54[20], i55[20], i56[20], i57[20],
i58[20], i59[20], i5A[20], i5B[20], i5C[20], i5D[20], i5E[20], i5F[20],
i60[20], i61[20], i62[20], i63[20], i64[20], i65[20], i66[20], i67[20],
i68[20], i69[20], i6A[20], i6B[20], i6C[20], i6D[20], i6E[20], i6F[20],
i70[20], i71[20], i72[20], i73[20], i74[20], i75[20], i76[20], i77[20],
i78[20], i79[20], i7A[20], i7B[20], i7C[20], i7D[20], i7E[20], i7F[20],
i80[20], i81[20], i82[20], i83[20], i84[20], i85[20], i86[20], i87[20],
i88[20], i89[20], i8A[20], i8B[20], i8C[20], i8D[20], i8E[20], i8F[20],
i90[20], i91[20], i92[20], i93[20], i94[20], i95[20], i96[20], i97[20],
i98[20], i99[20], i9A[20], i9B[20], i9C[20], i9D[20], i9E[20], i9F[20],
iA0[20], iA1[20], iA2[20], iA3[20], iA4[20], iA5[20], iA6[20], iA7[20],
iA8[20], iA9[20], iAA[20], iAB[20], iAC[20], iAD[20], iAE[20], iAF[20],
iB0[20], iB1[20], iB2[20], iB3[20], iB4[20], iB5[20], iB6[20], iB7[20],
iB8[20], iB9[20], iBA[20], iBB[20], iBC[20], iBD[20], iBE[20], iBF[20],
iC0[20], iC1[20], iC2[20], iC3[20], iC4[20], iC5[20], iC6[20], iC7[20],
iC8[20], iC9[20], iCA[20], iCB[20], iCC[20], iCD[20], iCE[20], iCF[20],
iD0[20], iD1[20], iD2[20], iD3[20], iD4[20], iD5[20], iD6[20], iD7[20],
iD8[20], iD9[20], iDA[20], iDB[20], iDC[20], iDD[20], iDE[20], iDF[20],
iE0[20], iE1[20], iE2[20], iE3[20], iE4[20], iE5[20], iE6[20], iE7[20],
iE8[20], iE9[20], iEA[20], iEB[20], iEC[20], iED[20], iEE[20], iEF[20],
iF0[20], iF1[20], iF2[20], iF3[20], iF4[20], iF5[20], iF6[20], iF7[20],
iF8[20], iF9[20], iFA[20], iFB[20], iFC[20], iFD[20], iFE[20], iFF[20]
}, S);
endmodule
/* VERY VERY BRAIN-UNFRIENDLY CODE ENDS*/
